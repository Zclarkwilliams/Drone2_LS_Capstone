`timescale 1ns / 1ns

/**
 * ECE 412-413 Capstone Winter/Spring 2018
 * Team 32 Drone2 SOC
 * Ethan Grinnell, Brett Creeley, Daniel Christiansen, Kirk Hooper, Zachary Clark-Williams
 */

/**
 * drone2 - Top level module for the drone controller.
 *
 * Outputs:
 * @motor_1_pwm: signal to drive the ESC connected to motor 1
 * @motor_2_pwm: signal to drive the ESC connected to motor 2
 * @motor_3_pwm: signal to drive the ESC connected to motor 3
 * @motor_4_pwm: signal to drive the ESC connected to motor 4
 *
 * Inputs:
 * @throttle_pwm: signal from throttle on the rc/receiver
 * @yaw_pwm: signal from yaw on the rc/receiver
 * @roll_pwm: signal from roll on the rc/receiver
 * @pitch_pwm: signal from pitch on the rc/receiver
 * @resetn: top level reset signal
 * @led_data_out: connects to the on board LEDs for the MachX03
 *
 * Inouts:
 * @sda: serial data line to the IMU
 * @scl: serial clock line to the IMU
 */

 `include "common_defines.v"

module drone2 (
	output wire motor_1_pwm,
	output wire motor_2_pwm,
	output wire motor_3_pwm,
	output wire motor_4_pwm,
	input wire throttle_pwm,
	input wire yaw_pwm,
	input wire roll_pwm,
	input wire pitch_pwm,
	input wire resetn,
	output wire rstn_imu,
	output wire [7:0]led_data_out,
	inout wire sda_1,
	inout wire sda_2,
	inout wire scl_1,
	inout wire scl_2);

	/* TODO: Figure out what these bit widths actually need to be
	 *		 and move them to the common_defines.v file.
	 */
	localparam REC_VAL_BIT_WIDTH = 8;   // values from receiver
	localparam PID_RATE_BIT_WIDTH = 16; // values from body frame controller
	localparam RATE_BIT_WIDTH = 16;     // values from angle controller
	localparam IMU_VAL_BIT_WIDTH = 16;  // values from IMU

	// values from receiver to angle_controller
	wire [REC_VAL_BIT_WIDTH-1:0] throttle_val;
	wire [REC_VAL_BIT_WIDTH-1:0] yaw_val;
	wire [REC_VAL_BIT_WIDTH-1:0] roll_val;
	wire [REC_VAL_BIT_WIDTH-1:0] pitch_val;

	// values from angle_controller to body_frame_controller
	wire [RATE_BIT_WIDTH-1:0] throttle_target_rate;
	wire [RATE_BIT_WIDTH-1:0] yaw_target_rate;
	wire [RATE_BIT_WIDTH-1:0] roll_target_rate;
	wire [RATE_BIT_WIDTH-1:0] pitch_target_rate;
	wire [RATE_BIT_WIDTH-1:0] roll_angle_error;
	wire [RATE_BIT_WIDTH-1:0] pitch_angle_error;

	// values from the IMU
	wire [IMU_VAL_BIT_WIDTH-1:0] x_linear_rate;
	wire [IMU_VAL_BIT_WIDTH-1:0] y_linear_rate;
	wire [IMU_VAL_BIT_WIDTH-1:0] z_linear_rate;
	wire [IMU_VAL_BIT_WIDTH-1:0] x_rotation;
	wire [IMU_VAL_BIT_WIDTH-1:0] y_rotation;
	wire [IMU_VAL_BIT_WIDTH-1:0] z_rotation;
	wire [IMU_VAL_BIT_WIDTH-1:0] x_rotation_rate;
	wire [IMU_VAL_BIT_WIDTH-1:0] y_rotation_rate;
	wire [IMU_VAL_BIT_WIDTH-1:0] z_rotation_rate;
	wire [IMU_VAL_BIT_WIDTH-1:0] x_linear_accel;
	wire [IMU_VAL_BIT_WIDTH-1:0] y_linear_accel;
	wire [IMU_VAL_BIT_WIDTH-1:0] z_linear_accel;

	// values from the body_frame_controller to the motor_mixer
	wire [PID_RATE_BIT_WIDTH-1:0] yaw_rate;
	wire [PID_RATE_BIT_WIDTH-1:0] roll_rate;
	wire [PID_RATE_BIT_WIDTH-1:0] pitch_rate;

	// values from motor_mixer to pwm_generator
	wire [`MOTOR_RATE_BIT_WIDTH-1:0] motor_1_rate;
	wire [`MOTOR_RATE_BIT_WIDTH-1:0] motor_2_rate;
	wire [`MOTOR_RATE_BIT_WIDTH-1:0] motor_3_rate;
	wire [`MOTOR_RATE_BIT_WIDTH-1:0] motor_4_rate;

	wire imu_good;
	wire iimu_data_valid;

	// status signals from angle_controller
	wire ac_valid_strobe;
	wire ac_active;

	// status signals from body_frame_controller
	wire bf_valid_strobe;
	wire bf_active;

	wire sys_clk;
	// TODO: Determine if we should stick with this clock rate (slower? faster?)
	defparam OSCH_inst.NOM_FREQ = "38.00";
	OSCH OSCH_inst (.STDBY(1'b0),
       			    .OSC(sys_clk),
       			    .SEDSTDBY());

	us_clk us_clk_divider (
		.us_clk(us_clk),
		.sys_clk(sys_clk),
		.resetn(resetn));


	bno055_driver	i(
		.scl_1(scl_1),                   //  I2C EFB SDA wires, Primary EFB
		.sda_1(sda_1),                   //  I2C EFB SDA wires, Primary EFB
		.scl_2(scl_2),                   //  I2C EFB SDA wires, Secondary EFB
		.sda_2(sda_2),                   //  I2C EFB SDA wires, Secondary EFB
		.rstn(resetn),                   //  async negative reset signal 0 = reset, 1 = not reset
		.led_data_out(led_data_out),     //  Module LED Status output -  //////////////////// Changed for testing, need to enable and feed LEDs somehow. /////////////////////
		.sys_clk(sys_clk),               //  master clock
		.rstn_imu(rstn_imu),             //  Low active reset signal to IMU hardware to trigger reset
		.imu_good(imu_good),             //  The IMU is either in an error or initial bootup states, measurements not yet active
		.imu_data_valid(imu_data_valid), //  Bit that indicates that the IMU data presented is valid, deasserted momentarily at 10ms polling interval and IMU burst read completion
		.gyro_rate_x(x_rotation_rate),   //  Rotation rate on X-Axis (Pitch rate)Precision: 1 Dps = 16 LSB
		.gyro_rate_y(y_rotation_rate),   //  Rotation rate on Y-Axis (Roll rate) Precision: 1 Dps = 16 LSB
		.gyro_rate_z(z_rotation_rate),   //  Rotation rate on Z-Axis (Yaw rate)  Precision: 1 Dps = 16 LSB
		.euler_angle_x(x_rotation),      //  Euler angle X-Axis       Pitch      Precision: 1 Deg = 16 LSB
		.euler_angle_y(y_rotation),      //  Euler angle Y-Axis       Roll       Precision: 1 Deg = 16 LSB
		.euler_angle_z(z_rotation),      //  Euler angle Z-Axis       Yaw        Precision: 1 Deg = 16 LSB
		.linear_accel_x(x_linear_accel), //  Linear Acceleration X-Axis          Precision: 1 m/s^2 = 100 LSB
		.linear_accel_y(y_linear_accel), //  Linear Acceleration Y-Axis          Precision: 1 m/s^2 = 100 LSB
		.linear_accel_z(z_linear_accel), //  Linear Acceleration Z-Axis          Precision: 1 m/s^2 = 100 LSB
		.x_velocity(x_linear_rate),
		.y_velocity(y_linear_rate),
		.z_velocity(z_linear_rate)
		);

	receiver receiver (
		.throttle_val(throttle_val),
		.yaw_val(yaw_val),
		.roll_val(roll_val),
		.pitch_val(pitch_val),
		.throttle_pwm(throttle_pwm),
		.yaw_pwm(yaw_pwm),
		.roll_pwm(roll_pwm),
		.pitch_pwm(pitch_pwm),
		.us_clk(us_clk),
		.resetn(resetn));

	angle_controller #(
		.RATE_BIT_WIDTH(RATE_BIT_WIDTH),
		.REC_VAL_BIT_WIDTH(REC_VAL_BIT_WIDTH),
		.IMU_VAL_BIT_WIDTH(IMU_VAL_BIT_WIDTH))
	angle_controller (
		.throttle_rate_out(throttle_target_rate),
		.yaw_rate_out(yaw_target_rate),
		.roll_rate_out(roll_target_rate),
		.pitch_rate_out(pitch_target_rate),
		.pitch_angle_error(pitch_angle_error),
		.roll_angle_error(roll_angle_error),
		.complete_signal(ac_valid_strobe),
		.active_signal(ac_active),
		.throttle_target(throttle_val),
		.yaw_target(yaw_val),
		.yaw_actual(x_rotation),
		.roll_target(roll_val),
		.pitch_target(pitch_val),
		.pitch_actual(x_rotation),
		.roll_actual(y_rotation),
		.resetn(resetn),
		.state(state),
		.start_signal(1'b1), // changed for testing, should be imu_data_valid
		.us_clk(us_clk));

/*
	body_frame_controller #(
		.PID_RATE_BIT_WIDTH(PID_RATE_BIT_WIDTH),
		.IMU_VAL_BIT_WIDTH(IMU_VAL_BIT_WIDTH),
		.PID_RATE_BIT_WIDTH(PID_RATE_BIT_WIDTH))
	body_frame_controller (
		.yaw_rate_out(yaw_rate),
		.roll_rate_out(roll_rate),
		.pitch_rate_out(pitch_rate),
		.complete_signal(bf_valid_strobe),
		.yaw_target(yaw_target_rate),
		.roll_target(roll_target_rate),
		.pitch_target(pitch_target_rate),
		.roll_rotation(x_rotation),
		.pitch_rotation(y_rotation),
		.yaw_rotation(z_rotation),
		.roll_angle_error(roll_angle_error),
		.pitch_angle_error(pitch_angle_error),
		.start_signal(ac_valid_strobe),
		.resetn(resetn),
		.us_clk(us_clk));
*/

	motor_mixer motor_mixer (
		.motor_1_rate(motor_1_rate),
		.motor_2_rate(motor_2_rate),
		.motor_3_rate(motor_3_rate),
		.motor_4_rate(motor_4_rate),
/*		// test connections
		.throttle_rate({4'h0, throttle_val, 4'h0}),
		.yaw_rate({4'h0, yaw_val, 4'h0}),
		.roll_rate({4'h0, roll_val, 4'h0}),
		.pitch_rate({4'h0, pitch_val, 4'h0}),
*/

		.throttle_rate(throttle_target_rate),
		.yaw_rate(yaw_target_rate),
		.roll_rate(roll_target_rate),
		.pitch_rate(pitch_target_rate),


		.sys_clk(sys_clk),
		.rst_n(resetn));

	// For now when in reset all LEDs are on
	//assign led_data_out = (!resetn) ? 8'h00 : 8'hFF;
	//assign led_data_out = ~throttle_target_rate[9:2];
	//assign led_data_out = {3'b111, ~state};
	//assign led_data_out = ~throttle_val;

	pwm_generator pwm_generator (
		.motor_1_pwm(motor_1_pwm),
		.motor_2_pwm(motor_2_pwm),
		.motor_3_pwm(motor_3_pwm),
		.motor_4_pwm(motor_4_pwm),
		.state_out(state_out),

		/*
		.motor_1_rate(throttle_val),
		.motor_2_rate(roll_val),
		.motor_3_rate(pitch_val),
		.motor_4_rate(yaw_val),
		*/

		.motor_1_rate(motor_1_rate),
		.motor_2_rate(motor_2_rate),
		.motor_3_rate(motor_3_rate),
		.motor_4_rate(motor_4_rate),


		.us_clk(us_clk),
		.resetn(resetn));

endmodule

