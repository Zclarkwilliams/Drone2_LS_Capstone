/**
 * ECE 412-413 Capstone Winter/Spring 2018
 * Team 32 Drone2 SOC
 * Ethan Grinnell, 
 * Brett Creeley, 
 * Daniel Christiansen, 
 * Kirk Hooper, 
 * Zachary Clark-Williams
 */
 
/**
 * Inputs:
 * (Target rates/angles are from the receiver module)
 * @throttle_target: 8-bit target rate from receiver module ranging from 0-250
 * @yaw_target: 8-bit target rate from receiver module ranging from 0-250
 * @pitch_target: 8-bit target angle from receiver module ranging from 0-250
 * @roll_target: 8-bit target angle from receiver module  ranging from 0-250
 * (Actual rates/angles are from the bno55_driver(IMU))
 * @yaw_actual: 16-bit, 2's complement fixed point [s11.4] actual rate in degrees
 * @pitch_actual: 16-bit, 2's complement fixed point [s11.4] actual rate in degrees
 * @roll_actual: 16-bit, 2's complement fixed point [s11.4] actual rate in degrees
 *
 * Outputs:
 * (Output rates are represented as 16-bit, 2's complement fixed point [s11.4])
 * @throttle_rate_out: limited to rate (>= 0) and represented as a scalar
 * @yaw_rate_out: limited yaw rate in degrees/second
 * @pitch_rate_out: limited pitch rate in degrees/second
 * @roll_rate_out: limited roll rate in degrees/second
 * (Output errors are represented as 16-bit, 2's complement fixed point [s11.4])
 * @pitch_angle_error: difference between the target and actual scaled
 * @roll_angle_error: difference between the target and actual scaled
 * (Signals used for module synchronization)
 * @complete_signal: Set high when the most recent calculation is done
 * @active_signal: Set high when currently calculating the next outputs
 * TODO:
 *		Clean up defines/localparams
 *		Rate limits???
 *		Optimize resource usage?
 */
`timescale 1ns / 1ns

`include "common_defines.v"

module angle_controller (
	output reg signed [`RATE_BIT_WIDTH-1:0] throttle_rate_out,
	output reg signed [`RATE_BIT_WIDTH-1:0] yaw_rate_out,
	output reg signed [`RATE_BIT_WIDTH-1:0] pitch_rate_out,
	output reg signed [`RATE_BIT_WIDTH-1:0] roll_rate_out,
	output reg signed [`RATE_BIT_WIDTH-1:0] pitch_angle_error,
	output reg signed [`RATE_BIT_WIDTH-1:0] roll_angle_error,
	output reg complete_signal,
	output reg active_signal,
	//output reg [4:0] state,
	input wire [`REC_VAL_BIT_WIDTH-1:0] throttle_target,
	input wire [`REC_VAL_BIT_WIDTH-1:0] yaw_target,
	input wire [`REC_VAL_BIT_WIDTH-1:0] pitch_target,
	input wire [`REC_VAL_BIT_WIDTH-1:0] roll_target,
	input wire signed [`RATE_BIT_WIDTH-1:0] yaw_actual /* synthesis syn_force_pads=1 syn_noprune=1*/ ,
	input wire signed [`RATE_BIT_WIDTH-1:0] pitch_actual,
	input wire signed [`RATE_BIT_WIDTH-1:0] roll_actual,
	input wire resetn,
	input wire start_signal,
	input wire us_clk);

	// TODO: Use decimal values instead to avoid having to comment
	// rate limits (16-bit, 2's complement, 12-bit integer, 4-bit fractional)
	localparam signed
		THROTTLE_MAX = 16'h0fa0, // 250
		YAW_MAX =      16'h0640, // 100
		YAW_MIN =      16'hf9C0, // -100
		PITCH_MAX =    16'h0640, // 100
		PITCH_MIN =    16'hf9C0, // -100
		ROLL_MAX =     16'h0640, // 100
		ROLL_MIN =     16'hf9C0; // -100

	// scale factors (16-bit, 2's complement, 12-bit integer, 4-bit fractional)
	localparam signed
		THROTTLE_SCALE = 16'd1,
		YAW_SCALE =      16'd48,
		ROLL_SCALE =     16'd32,
		PITCH_SCALE =    16'd32;

	// TODO: Remove unused variables
	// working registers
	reg signed [`RATE_BIT_WIDTH-1:0] mapped_throttle, mapped_yaw, mapped_roll, mapped_pitch;
	reg signed [`RATE_BIT_WIDTH-1:0] new_mapped_throttle, new_mapped_yaw, new_mapped_roll, new_mapped_pitch;
	reg signed [`RATE_BIT_WIDTH-1:0] scaled_throttle, scaled_yaw, scaled_roll, scaled_pitch;
	reg signed [`REC_VAL_BIT_WIDTH-1:0] latched_throttle, latched_yaw, latched_pitch, latched_roll;


	// state names
	localparam
		STATE_WAITING =  5'b00001,
		STATE_MAPPING =  5'b00010,
		STATE_SCALING =  5'b00100,
		STATE_LIMITING = 5'b01000,
		STATE_COMPLETE = 5'b10000;

	// state variables
	reg [4:0] state, next_state;

	reg start_flag = 1'b0;

	// latch start signal
	always @(posedge us_clk or negedge resetn) begin
		if(!resetn)
			start_flag <= 1'b0;
		else if(start_signal && !start_flag)
			start_flag <= 1'b1;
		else if(!start_signal && start_flag) begin
			if(state != STATE_WAITING) begin
				start_flag <= 1'b0;
			end
		end
		else
			start_flag <= start_flag;
	end

	// update state
	always @(posedge us_clk or negedge resetn) begin
		if(!resetn) begin
			state <= STATE_WAITING;
			latched_throttle <= 16'h0000;
			latched_yaw <= 16'h00000;
			latched_pitch <= 16'h0000;
			latched_roll <= 16'h0000;
		end
		else begin
			state <= next_state;
			latched_throttle <= throttle_target;
			latched_yaw <= yaw_target;
			latched_pitch <= pitch_target;
			latched_roll <= roll_target;

		end

	end

	// next state logic
	always @(*) begin
		case(state)
			STATE_WAITING: begin
				if(start_flag)
					next_state = STATE_MAPPING;
				else
					next_state = STATE_WAITING;
			end
			STATE_MAPPING: begin
				next_state = STATE_SCALING;
			end
			STATE_SCALING: begin
				next_state = STATE_LIMITING;
			end
			STATE_LIMITING: begin
				next_state = STATE_COMPLETE;
			end
			STATE_COMPLETE: begin
				next_state = STATE_WAITING;
			end
			default: begin
				next_state = STATE_WAITING;
			end
		endcase
	end



	// output logic
	always @(posedge us_clk or negedge resetn) begin
		if(!resetn) begin
			// reset values
			yaw_rate_out <= 16'h0000;
			roll_rate_out <= 16'h0000;
			pitch_rate_out <= 16'h0000;

		end
		else begin
			case(state)
				STATE_WAITING: begin
					complete_signal <= 1'b0;
					active_signal <= 1'b0;
				end
				STATE_MAPPING: begin
					complete_signal <= 1'b0;
					active_signal <= 1'b1;

					mapped_throttle <= {4'h0, latched_throttle, 4'h0};
					// input values mapped from 0 - 250 to -31.25 - 31.25
					mapped_yaw <= $signed({6'b0, latched_yaw, 2'b0}) - $signed(16'd500);
					// roll value from IMU is flipped, add instead of subtract (do this in bfc too?)
					mapped_roll <= ($signed({6'b0, latched_roll, 2'b0}) - $signed(16'd500)) + $signed(roll_actual);
					mapped_pitch <= ($signed({6'b0, latched_pitch, 2'b0}) - $signed(16'd500)) - $signed(pitch_actual);
				end
				STATE_SCALING: begin
					complete_signal <= 1'b0;
					active_signal <= 1'b1;

					// the decimal point should be shifted...
					scaled_throttle <= (mapped_throttle * THROTTLE_SCALE);
					scaled_yaw <= (mapped_yaw * YAW_SCALE) >>> 4;
					scaled_roll <= (mapped_roll * ROLL_SCALE) >>> 4;
					scaled_pitch <= (mapped_pitch * PITCH_SCALE) >>> 4;
				end
				STATE_LIMITING: begin
					complete_signal <= 1'b0;
					active_signal <= 1'b1;

					//TODO: Add throttle min checking
					// apply rate limits
					if(scaled_throttle > THROTTLE_MAX)
						throttle_rate_out <= THROTTLE_MAX;
					else
						throttle_rate_out <= scaled_throttle;

					if(scaled_yaw > YAW_MAX)
						yaw_rate_out <= YAW_MAX;
					else if(scaled_yaw < YAW_MIN)
						yaw_rate_out <= YAW_MIN;
					else
						yaw_rate_out <= scaled_yaw;

					if(scaled_roll > ROLL_MAX)
						roll_rate_out <= ROLL_MAX;
					else if(scaled_roll < ROLL_MIN)
						roll_rate_out <= ROLL_MIN;
					else
						roll_rate_out <= scaled_roll;

					if(scaled_pitch > PITCH_MAX)
						pitch_rate_out <= PITCH_MAX;
					else if(scaled_pitch < PITCH_MIN)
						pitch_rate_out <= PITCH_MIN;
					else
						pitch_rate_out <= scaled_pitch;

					pitch_angle_error <= mapped_pitch;
					roll_angle_error <= mapped_roll;
				end
				STATE_COMPLETE: begin
					complete_signal <= 1'b1;
					active_signal <= 1'b0;
				end
				default: begin
					pitch_rate_out <= 16'h0000;
					yaw_rate_out <= 16'h0000;
					roll_rate_out <= 16'h0000;
					throttle_rate_out <= 16'h0000;
				end
			endcase
		end
	end

endmodule

